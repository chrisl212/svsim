module prop;

  assert property ((in & in_2) |-> 2) begin

  end

endmodule
